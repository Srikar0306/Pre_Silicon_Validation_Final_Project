package fifo_pkg;

	`include "async_seq_item.sv"
`include "async_sequence_basetest.sv"

	`include "async_sequencer.sv"
	`include "async_driver.sv"
	`include "write_monitor.sv"
	`include "read_monitor.sv"
	`include "async_write_agent.sv"
	`include "async_read_agent.sv"
	`include "async_scoreboard.sv"

		
endpackage
